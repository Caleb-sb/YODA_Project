//------------------------------------------------------------------------------
// File name	:	top.v
// Module Name	:	top
// Function		:	Implements FSM to output arpeggio or just base note
// Coder		:	Caleb Bredekamp [BRDCAL003]
// Comments		:	Adapted from template given by Keegan Crankshaw:
//					https://github.com/UCT-EE-OCW/EEE4120F-Pracs
//------------------------------------------------------------------------------
module SD_Controller(

	);
endmodule